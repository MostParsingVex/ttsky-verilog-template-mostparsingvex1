/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_mostparsingvex1(
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  wire rst;
  assign rst = !rst_n;
  wire[7:0] data_in;
  //assign data_in[3:0] = ui_in[3:0];
  //assign data_in[7:4] = 4'h0;
  assign data_in[4:0] = ui_in[4:0]
  assign data_in[7:5] = 3'h0;
  amx_core1 U0( .clk( clk ), .rst( rst ), .data_in( data_in ), .data_out( uo_out ) );

  // All output pins must be assigned. If not used, assign to 0.
  //assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = ui_in | uio_in;
  assign uio_oe = 8'hff;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};

endmodule
